`timescale 1ns/1ns

module glbl_sink ();

    wire rst;

    assign rst = glbl.rst;

endmodule