-- Invalid VHDL file

invalid_statement;
