

module test_parameters #(
    parameter WIDTH_IN = 8,
    parameter WIDTH_OUT = 8
) (
    input  [WIDTH_IN-1:0]   IN,
    output [WIDTH_OUT-1:0]  OUT
);

endmodule
